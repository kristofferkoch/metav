module mem;
   reg [7:0] bytes [255:0], shadow [255:0], single;
endmodule // mem
